* Monte Carlo simulation in NGSpice (Transient)
Vin in 0 DC 10V
R1 in out {R1}
R2 out 0 {R2}

* Define parameterized resistor values with Gaussian variation
.param mc_run = 0
.param R1 = 1k * (1 + gauss(0, 0.05))   ; 5% variation
.param R2 = 1k * (1 + gauss(0, 0.05))   ; 5% variation

* Transient analysis setup (simulate for 1ms)
.tran 0.1ms 1ms

.control
set filetype=ascii
destroy all
reset
* Create the output file for saving results
outf=open monte_output.txt

foreach i 1 100
  alterparam mc_run = $i
  run
  * Save output voltage to the file
  print v(out) > outf
end

* Close the output file
close outf
.endc

.end
